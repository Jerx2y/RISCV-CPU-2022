// execution
module EX (
    
);
    
endmodule