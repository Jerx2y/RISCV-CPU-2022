// Issue
`include "defines.v"

module Issue (
    input wire clk, rst, rdy

    // IFetcher
);



endmodule