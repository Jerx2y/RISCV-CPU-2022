// register module
module REG (
    
);
    
endmodule