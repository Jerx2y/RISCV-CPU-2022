// load store buffer
module LSB (
    
);
    
endmodule