// instruction fetch
module IF (
    
);
    
endmodule