// reorder buffer
module ROB (
    
);
    
endmodule