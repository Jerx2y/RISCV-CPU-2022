// instruction cache
module IC (
    
);
    
endmodule