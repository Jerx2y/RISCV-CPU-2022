// memory controller
module MC (
    
);
    
endmodule