// Decoder
module DC (
    
);



endmodule