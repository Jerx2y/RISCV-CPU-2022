// data cache
module DC (
    
);
    
endmodule