// instruction cache

module ICache (
    
);
    
endmodule