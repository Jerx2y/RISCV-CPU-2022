`include "defines.v"

module IFetch (
    input wire clk, rst, rdy,
    
    // Decoder
    

    // ICache
    input wire [31 : 0] ins,
);

reg [31 : 0] imm;

reg [31 : 0] pc;

always @(*) begin
    
end



endmodule