// reservation station
module RS (
    
);
    
endmodule